module tb_riscV();

endmodule
