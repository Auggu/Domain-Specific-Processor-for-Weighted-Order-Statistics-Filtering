module instr_rom #(
    parameter SIZE = 512
) (
    input i_clk,
    input i_rst,
    input [31:0] i_addr,
    output [31:0] o_out
);
endmodule

